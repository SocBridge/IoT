//jayaram
module test;
  initial
    begin
	$display("Welcome to SocBridge Semiconductors Pvt Ltd");
	$display("Bangalore");
    end

enmodule 
